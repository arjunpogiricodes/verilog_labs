


module random_counter(clk,reset,count);

// declaration of ports
