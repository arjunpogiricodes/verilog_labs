


module fsm_code_style_4(clk,reset,d_in,d_out);

// declaring the input and output ports

  input clk,reset,d_in;
  output d_out;
// parameter and regs declaration

   parameter s0=3'b000,s1=3'b100,s2=
